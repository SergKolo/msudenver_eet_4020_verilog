module veriogAND(Fv,Av,Bv);
    input Av,Bv;
	 output Fv;
	 and v_and(Fv,Av,Bv);
endmodule
